library ieee;
use ieee.numeric_bit.all;

entity ula1bit is
    port (
        a         : in bit;
        b         : in bit;
        cin       : in bit;
        ainvert   : in bit;
        binvert   : in bit;
        operation : in bit_vector(1 downto 0);
        result    : out bit;
        cout      : out bit;
        overflow  : out bit
    );
end entity ula1bit;

architecture structural of ula1bit is
    -- Internal signals inputs (invert or not)
    signal a_val, b_val : bit;
    
    -- Results from sub-blocks
    signal res_and : bit;
    signal res_or  : bit;
    signal res_add : bit; -- Sum from adder
    signal c_out_s : bit; -- Carry out from adder

begin
    -- Input Inversion Logic (Multiplexers)
    -- If ainvert=1, use NOT a; else use a.
    a_val <= not a when ainvert = '1' else a;
    b_val <= not b when binvert = '1' else b;

    -- Logic Operations
    res_and <= a_val and b_val;
    res_or  <= a_val or b_val;

    -- Arithmetic Operation (Full Adder Instantiation)
    adder: entity work.fulladder
        port map (
            a    => a_val,
            b    => b_val,
            cin  => cin,
            s    => res_add,
            cout => c_out_s
        );

    -- Output Multiplexer (Selects result based on 'operation')
    -- 00: AND
    -- 01: OR
    -- 10: ADD
    -- 11: Pass B (Passes the processed B value)
    with operation select result <=
        res_and when "00",
        res_or  when "01",
        res_add when "10",
        b       when "11"; -- Pass B

    -- Carry Out is generated by the adder
    cout <= c_out_s;

    -- Overflow Detection
    -- For the MSB, overflow occurs if Carry In != Carry Out
    overflow <= cin xor c_out_s;

end architecture structural;